library IEEE;
	use IEEE.std_logic_1164.ALL;
	use IEEE.std_logic_arith.ALL;
	use IEEE.std_logic_unsigned.ALL;

library hdl_library_CommonFunctions;
	use hdl_library_CommonFunctions.MathHelpers.all;

library hdl_library_ClockGenerator;
	use hdl_library_ClockGenerator.all;


library hdl_library_DSP_Filter_FIR;
	use hdl_library_DSP_Filter_FIR.all;

entity FIR_CoreTB is
end entity; --FIR_CoreTB

architecture arch of FIR_CoreTB is

	constant G_CLOCK_FREQUENCY 					: integer := 100E6;

	constant C_FIR_FILTER_ORDER 				: integer := 16;

	constant C_DATA_IN_WIDTH 					: integer := 32;
	constant C_DATA_OUT_WIDTH 					: integer := 32;

	constant C_COEFF_WIDTH 						: integer := 32;


	signal clock 								: std_logic := '0';
	signal clock_n 								: std_logic := '0';
	signal enable 								: std_logic := '0';

	type T_COEFF_ROM is array(0 to C_FIR_FILTER_ORDER - 1) of std_logic_vector(C_COEFF_WIDTH - 1 downto 0);
	signal coeff_ROM 							: T_COEFF_ROM := (others => (others => '0'));

	signal xn 									: std_logic_vector(C_DATA_IN_WIDTH - 1 downto 0) := (others => '0');
	signal xn_nd 								: std_logic := '0';
	
	signal yn 									: std_logic_vector(C_DATA_OUT_WIDTH - 1 downto 0) := (others => '0');
	signal yn_valid 							: std_logic := '0';

	signal current_coefficient 					: std_logic_vector(C_COEFF_WIDTH - 1 downto 0) := (others => '0');
	signal current_coefficient_address 			: std_logic_vector(log2(C_FIR_FILTER_ORDER) - 1 downto 0) := (others => '0');

begin

	clock <= not clock after (1 sec / G_CLOCK_FREQUENCY) / 2;
	clock_n <= not clock;

	enable <= '1' after 100 ns;

	dut : entity hdl_library_DSP_Filter_FIR.FIR_Core
	generic map
	(
		C_FIR_FILTER_ORDER 					=> C_FIR_FILTER_ORDER,

		C_DATA_IN_WIDTH 					=> C_DATA_IN_WIDTH,
		C_DATA_OUT_WIDTH 					=> C_DATA_OUT_WIDTH,

		C_COEFF_WIDTH 						=> C_COEFF_WIDTH
	)
	port map
	(
		clock 								=> clock,
		enable 								=> enable,

		xn 									=> xn,
		xn_nd 								=> xn_nd,

		yn 									=> yn,
		yn_valid 							=> yn_valid,

		current_coefficient 				=> current_coefficient,
		current_coefficient_address 		=> current_coefficient_address


		--ready 								=> ready
	);

end architecture; -- arch